	module Mem(Clk,BE,CS,RW,Addr,DataIn,Reset,DataOut,DataReady);
	input        Clk,CS,RW,Reset;
	input[3:0]   BE;
	input[31:2]  Addr;
	input[31:0]  DataIn;
	output[31:0] DataOut;
	output       DataReady;
	
	(*ram_init_file = "D:\new\Mem.mif"*)
	reg[31:0]    memory[31:0];
	reg[31:0]    DataOut;
	
	assign DataReady=1;
	
	always@(posedge Clk or posedge Reset)
	  if(Reset)begin
	    memory[0]<=32'b00000000000000000000000000000000;
	    memory[1]<=32'b00000000000000000000000000000000;
	    memory[2]<=32'b00000000000000000000000000000000;
	    memory[3]<=32'b00000000000000000000000000000000;
	    memory[4]<=32'b00000000000000000000000000000000;
	    memory[5]<=32'b00000000000000000000000000000000;
	    memory[6]<=32'b00000000000000000000000000000000;
	    memory[7]<=32'b00111100000010001011111111000000;
	    memory[8]<=32'b00111100000100000000000000000110;
	    memory[9]<=32'b00111100000100010000000000000100;
	   memory[10]<=32'b00111100000100100000000000000001;
	   memory[11]<=32'b00111100000101010000000000000000;
	   memory[12]<=32'b00000010000100001001000000100110;
	   memory[13]<=32'b00000010011100001000000000001011;
	   memory[14]<=32'b00100110100101000000000000000100;
	   memory[15]<=32'b00000001000010001010000000100001;
	   memory[16]<=32'b10001101000101010000000000000000;
	   memory[17]<=32'b10001101000101100000000000000100;
	   memory[18]<=32'b00000001001101011011000000100011;
	   memory[19]<=32'b00011101001000000000000000000100;
	   memory[20]<=32'b00000010111010101000000000001011;
	   memory[21]<=32'b00000010101101101000000000001011;
	   memory[22]<=32'b00000010110101111000000000001011;
	   memory[23]<=32'b10101101000101010000000000000000;
	   memory[24]<=32'b10101101000101100000000000000100;
	   memory[25]<=32'b00000001000010001010000000100011;
	   memory[26]<=32'b00000010011100111001000000100011;
	   memory[27]<=32'b00011010011000000000000000000010;
	   memory[28]<=32'b00001011111100000000000000100111;
	   memory[29]<=32'b00000010000100001001000000100011;
	   memory[30]<=32'b00011010000000000000000000000010;
	   memory[31]<=32'b00001011111100000000000000101010;
	  end
	  else if(Clk)
	  begin
	    if(RW)begin
	      memory[Addr[6:2]][31:16]<=(BE[3:2]==2'b11)?DataIn[31:16]:16'b0;
	      memory[Addr[6:2]][15:8] <=(BE[1]==1'b1)?DataIn[15:8]:8'b0;
	      memory[Addr[6:2]][7:0] <=DataIn[7:0];
	    end
	    else begin
	      DataOut[31:16]<=(BE[3:2]==2'b11)?memory[Addr[6:2]][31:16]:16'b0;
	      DataOut[15:8] <=(BE[1]==1'b1)?memory[Addr[6:2]][15:8]:8'b0;
	      DataOut[7:0]  <=memory[Addr[6:2]][7:0];
	    end
	  end
	endmodule