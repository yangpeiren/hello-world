//8λ�첽����ͨ�Ž�����
//��ģ�鰴�չ̶��Ĳ����ʣ�9600*16bit/s�������մ����źţ�
//������ֹʽ�첽Э�飬��ʼλΪһλ�ĵ͵�ƽ�����ݳ���Ϊ8λ����������żУ��λ��ֹͣλΪ2λ�ߵ�ƽ��
//�����ɺ���������źţ��Լ�������ݣ�
module rs_232_in(clk, shiftin, in_data, data_finish);

	input clk;					//����ʱ�ӣ�(9600*16)hz
	input shiftin;				//�������������

	output[7:0] in_data;		//��������ź�8λ�������
	output data_finish;			//���ݽ��ܽ����ź�
	
	reg[7:0] in_data;			//�������ݼĴ���
	reg data_finish;			//���ݽ��ܽ����ź�
	reg flag;					//���ݽ���״̬�Ĵ�����0���ȴ�״̬��1������״̬��
	reg[7:0] count;				//���������

	always @(posedge clk)
	begin
		//�����������ڵȴ�״̬ʱ�����յ���ʼλ��?�źţ���״̬�Ĵ���Ϊ1���������״̬��
		if(flag == 0 && shiftin == 0)
			flag <= 1;
		//�����������ڽ���״̬ʱ,��������ʼ������
		else if(flag == 1)
			count <= count + 8'b1;
		//�����ź�λ��0��
		data_finish <= 0;
		//���ݽ����߼����֣�
		if((count[7:4] <= 8) && (count[3:0] == 0) && (flag == 1))  	//������������16��ʱ����ʼ�������ݣ�һ������8λ��
		begin
			in_data <= in_data >> 1;								//�Ĵ�����1λ��ѭ������	
			in_data[7] <= shiftin;								//�����յ�������д��Ĵ�����λ
		end
		else if((count[7:4] == 11) && (count[3:0] == 0))			//��������
		begin
			flag <= 0;											//�������ɽ���״̬����ȴ�״̬
			data_finish <= 1;									//������ܽ����ź�
			count <= 0;										//��������0
		end
	end
endmodule



