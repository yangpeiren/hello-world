module Constant(const4,const14,const31);
output[4:0] const14,const31;
output[31:0] const4;

assign const14=5'd14;
assign const31=5'd31;
assign const4 =32'd4;

endmodule
